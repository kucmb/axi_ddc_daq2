`timescale 1 ns / 1 ps

module ddc_quad(
    input clk,

    // assuming [29:16] Q, [13:0] I
    input [31:0] data_in_0,
    input [31:0] data_in_1,
    input [31:0] data_in_2,
    input [31:0] data_in_3,

    input [19:0] pinc,
    input [19:0] poff,
    input p_valid,

    output valid_out,
    output [63:0] data_out
);

    localparam LATENCY_P = 3;
    localparam LATENCY_SUM = 6;

    wire valid_in_dds;
    wire valid_out_ddc;

    wire [19:0] poff_0;
    wire [19:0] poff_1;
    wire [19:0] poff_2;
    wire [19:0] poff_3;

    wire [63:0] ddc_out_0;
    wire [63:0] ddc_out_1;
    wire [63:0] ddc_out_2;
    wire [63:0] ddc_out_3;

    wire [19:0] pinc_x2;
    wire [19:0] pinc_x3;
    wire [19:0] pinc_x4;

    // Valid signal management
    reg [LATENCY_P-1:0] p_valid_buf;
    reg [LATENCY_SUM-1:0] valid_out_buf;

    // Sum
    wire [29:0] i_03;
    wire [29:0] q_03;
    wire [29:0] i_12;
    wire [29:0] q_12;
    wire [30:0] i_tot;
    wire [30:0] q_tot;

    assign data_out = {q_tot[30], q_tot, i_tot[30], i_tot};

    always @(posedge clk) begin
        p_valid_buf = {p_valid_buf[LATENCY_P-2:0], p_valid};
    end
    assign valid_in_dds = p_valid_buf[LATENCY_P-1];

    always @(posedge clk) begin
        valid_out_buf = {valid_out_buf[LATENCY_SUM-2:0], valid_out_ddc};
    end
    assign valid_out = valid_out_buf[LATENCY_SUM-1];

    // Phase increment and offset calculation for quad-mode operation
    assign pinc_x4 = {pinc[17:0], 2'b0};
    assign pinc_x2 = {pinc[18:0], 1'b0};
    assign pinc_x3 = pinc + pinc_x2;
    
    // phase adder
    adder_phase add_0(
        .clk(clk),
        .a(poff),
        .b(20'b0),
        .s(poff_0)
    );

    adder_phase add_1(
        .clk(clk),
        .a(poff),
        .b(pinc),
        .s(poff_1)
    );

    adder_phase add_2(
        .clk(clk),
        .a(poff),
        .b(pinc_x2),
        .s(poff_2)
    );

    adder_phase add_3(
        .clk(clk),
        .a(poff),
        .b(pinc_x3),
        .s(poff_3)
    );

    // DDC instantiation
    ddc_core ddc_0(
        .clk(clk),
        .data_in(data_in_0),
        .valid_in(valid_in_dds),
        .phase_in({4'b0, poff_0, 4'b0, pinc_x4}),
        .valid_out(valid_out_ddc),
        .ddc_out(ddc_out_0)
    );

    ddc_core ddc_1(
        .clk(clk),
        .data_in(data_in_1),
        .valid_in(valid_in_dds),
        .phase_in({4'b0, poff_1, 4'b0, pinc_x4}),
        .ddc_out(ddc_out_1)
    );

    ddc_core ddc_2(
        .clk(clk),
        .data_in(data_in_2),
        .valid_in(valid_in_dds),
        .phase_in({4'b0, poff_2, 4'b0, pinc_x4}),
        .ddc_out(ddc_out_2)
    );

    ddc_core ddc_3(
        .clk(clk),
        .data_in(data_in_3),
        .valid_in(valid_in_dds),
        .phase_in({4'b0, poff_3, 4'b0, pinc_x4}),
        .ddc_out(ddc_out_3)
    );


    // Output adder
    adder_1st add_i_03(
        .clk(clk),
        .a(ddc_out_0[28:0]),
        .b(ddc_out_3[28:0]),
        .s(i_03)
    );

    adder_1st add_q_03(
        .clk(clk),
        .a(ddc_out_0[60:32]),
        .b(ddc_out_3[60:32]),
        .s(q_03)
    );

    adder_1st add_i_12(
        .clk(clk),
        .a(ddc_out_1[28:0]),
        .b(ddc_out_2[28:0]),
        .s(i_12)
    );

    adder_1st add_q_12(
        .clk(clk),
        .a(ddc_out_1[60:32]),
        .b(ddc_out_2[60:32]),
        .s(q_12)
    );

    adder_2nd add_i_tot(
        .clk(clk),
        .a(i_03),
        .b(i_12),
        .s(i_tot)
    );

    adder_2nd add_q_tot(
        .clk(clk),
        .a(q_03),
        .b(q_12),
        .s(q_tot)
    );

endmodule
